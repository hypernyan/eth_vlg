module tcp_vlg_rx 
  import
    ipv4_vlg_pkg::*,
    mac_vlg_pkg::*,
    tcp_vlg_pkg::*,
    eth_vlg_pkg::*;
(
  input logic clk,
  input logic rst,
  ipv4.in_rx  ipv4,
  tcp.out_rx  tcp
);
  enum logic [4:0] {idle_s, hdr_s, opt_s, pld_s, rst_s} fsm;

  logic fsm_rst;
  logic  [$clog2(TCP_HDR_LEN)+4:0] byte_cnt; // maximum 
  
  logic [tcp_vlg_pkg::TCP_HDR_LEN-1:0][7:0] hdr;
  logic [tcp_vlg_pkg::TCP_MAX_OPT_LEN-1:0][7:0] opt;

  logic [5:0] offset;
    // Latch header
  logic rst_reg;
  tcp_opt_field_t opt_field;
  tcp_opt_type_t cur_opt;

  length_t len, pld_byte_cnt;

  logic [7:0] opt_byte_cnt, opt_len;

  assign fsm_rst = rst || rst_reg;

  // TCP receive FSM
  // The state machine here is responsible for receiving TCP packets and parsing header and options
  // Main (20 bytes) header is generated by a simple shiftreg that triggers output when byte count reaches 20.
  // After the main header was latched, the FSM processes options if there are any (IHL > 5)
  // The options are specifissssssssssssed, so the FSM follows those specs
  // A present
  always_ff @ (posedge clk) begin
    if (fsm_rst) begin
      fsm          <= idle_s;
      byte_cnt     <= 0;
      pld_byte_cnt <= 0;
      tcp.strm     <= 0;
      tcp.meta     <= 0;
      offset       <= 0;
      opt_len      <= 0;
      cur_opt      <= tcp_opt_nop;
      opt_field    <= tcp_opt_field_kind;
      hdr          <= 0;
      rst_reg      <= 0;
      len          <= 0;
    end
    else begin
      hdr[tcp_vlg_pkg::TCP_HDR_LEN-1:1] <= hdr[tcp_vlg_pkg::TCP_HDR_LEN-2:0];
      hdr[0] <= ipv4.strm.dat;
      opt[tcp_vlg_pkg::TCP_MAX_OPT_LEN-1:1] <= opt[tcp_vlg_pkg::TCP_MAX_OPT_LEN-2:0];
      opt[0] <= ipv4.strm.dat;
            
      case (fsm)
        idle_s : begin
          if (ipv4.strm.val && ipv4.strm.sof && (ipv4.meta.ipv4_hdr.proto == TCP)) begin
            tcp.meta.mac_hdr  <= ipv4.meta.mac_hdr;
            tcp.meta.ipv4_hdr <= ipv4.meta.ipv4_hdr;
            len <= ipv4.meta.pld_len;
            fsm <= hdr_s;
          end    
        end
        hdr_s : begin
          byte_cnt <= byte_cnt + 1;
          if (byte_cnt == tcp_vlg_pkg::HDR_OPTIONS_POS-1) offset <= ipv4.strm.dat[7:4] << 2; // TCP offset field will be exactly at [7:4]. multiply by 4
          tcp.meta.pld_len <= len - offset; // calculate TCP payload length
          // choose the way to proceed based on offset and payload length:
          // - if offset is more then 5, there are TCP options, parse them
          // - if payload length is zero, reset the FSM
          // - if payload length is non-zero, process the payload
          if (byte_cnt == TCP_HDR_LEN - 2) begin
            fsm <= (offset == TCP_HDR_LEN) ? (tcp.meta.pld_len == 0) ? rst_s : pld_s : opt_s; 
            tcp.meta.tcp_hdr <= {hdr[18:0], ipv4.strm.dat};
          end
        end
        opt_s : begin
          byte_cnt <= byte_cnt + 1;
          // If there is no payload, skip it and process to reset state
          if (byte_cnt == offset - 2) fsm <= (tcp.meta.pld_len == 0) ? rst_s : pld_s;
          case (opt_field)
            tcp_opt_field_kind : begin
              case (ipv4.strm.dat)
                TCP_OPT_END : begin
                //  $display("Option kind: end");
                  opt_field <= tcp_opt_field_kind;
                  cur_opt <= tcp_opt_end;
                end
                TCP_OPT_NOP : begin
                //  $display("Option kind: NOP");
                  opt_field <= tcp_opt_field_kind;
                  cur_opt <= tcp_opt_nop;
                end
                TCP_OPT_MSS : begin
                //  $display("Option kind: MSS");
                  tcp.meta.tcp_opt.tcp_opt_pres.mss_pres <= 1;
                  opt_field <= tcp_opt_field_len;
                  cur_opt <= tcp_opt_mss;
                end
                TCP_OPT_WIN : begin
                //  $display("Option kind: wnd");
                  tcp.meta.tcp_opt.tcp_opt_pres.wnd_pres <= 1;
                  opt_field <= tcp_opt_field_len;
                  cur_opt <= tcp_opt_wnd; 
                end
                TCP_OPT_SACK_PERM : begin
                //  $display("Option kind: SACK Permitted");
                  tcp.meta.tcp_opt.tcp_opt_pres.sack_perm_pres <= 1;
                  opt_field <= tcp_opt_field_len;
                  cur_opt <= tcp_opt_sack_perm;
                end
                TCP_OPT_SACK : begin
                //  $display("Option kind: SACK");
                  tcp.meta.tcp_opt.tcp_opt_pres.sack_pres <= 1;
                  opt_field <= tcp_opt_field_len;
                  cur_opt <= tcp_opt_sack;  
                end
                TCP_OPT_TIMESTAMP : begin
                //  $display("Option kind: timestamp");
                  tcp.meta.tcp_opt.tcp_opt_pres.timestamp_pres <= 1;
                  opt_field <= tcp_opt_field_len;
                  cur_opt <= tcp_opt_timestamp;
                end
                default : begin
                  opt_field <= tcp_opt_field_kind;
                end
              endcase
              opt_byte_cnt <= 0;
            end
            tcp_opt_field_len : begin
              case (ipv4.strm.dat) // Only SACK has variable length
                10      : tcp.meta.tcp_opt.tcp_opt_sack.block_pres <= 4'b1000;
                18      : tcp.meta.tcp_opt.tcp_opt_sack.block_pres <= 4'b1100;
                26      : tcp.meta.tcp_opt.tcp_opt_sack.block_pres <= 4'b1110;
                34      : tcp.meta.tcp_opt.tcp_opt_sack.block_pres <= 4'b1111;
                default : tcp.meta.tcp_opt.tcp_opt_sack.block_pres <= 4'b0000;
              endcase
              opt_len <= ipv4.strm.dat - 2; // exclude kind and length bytes
              opt_field <= (ipv4.strm.dat == 2) ? tcp_opt_field_kind : tcp_opt_field_data;
            end
            tcp_opt_field_data : begin
              opt_byte_cnt <= opt_byte_cnt + 1;
              if (opt_byte_cnt == opt_len - 1) begin
                opt_field <= tcp_opt_field_kind;
                case (cur_opt)
                  tcp_opt_mss : begin
                  //  $display("MSS Option value: %d", opt_data[1:0]);
                    tcp.meta.tcp_opt.tcp_opt_mss.mss <= {opt[0], ipv4.strm.dat};
                  end
                  tcp_opt_wnd : begin
                  //  $display("Window Option value: %d", opt_data[0]);
                    tcp.meta.tcp_opt.tcp_opt_wnd.wnd <= ipv4.strm.dat;
                  end
                  tcp_opt_sack : begin
                      tcp.meta.tcp_opt.tcp_opt_sack.block[0] <= {opt[6:0], ipv4.strm.dat};
                    if (opt_byte_cnt == 6 || opt_byte_cnt == 14 || opt_byte_cnt == 22 || opt_byte_cnt == 30) begin
                      tcp.meta.tcp_opt.tcp_opt_sack.block[1:3]     <= tcp.meta.tcp_opt.tcp_opt_sack.block[0:2];
                    end
                  //  $display("SACK Option value: Begin: %h, End: %h", opt_data[7:4], opt_data[3:0]);
                  end
                  tcp_opt_timestamp : begin
                   // tcp.meta.tcp_opt.tcp_opt_timestamp.timestamp <= {hdr[0], ipv4.strm.dat};
                  end
                endcase
              end
            end
          endcase
        end
        pld_s : begin
          tcp.meta.pkt_start <= tcp.meta.tcp_hdr.tcp_seq_num;
          tcp.meta.pkt_stop  <= tcp.meta.tcp_hdr.tcp_seq_num + tcp.meta.pld_len;
          pld_byte_cnt <= pld_byte_cnt + 1;
          if (pld_byte_cnt == tcp.meta.pld_len - 1) fsm <= rst_s;
          tcp.meta.val <= 1;
          tcp.strm.dat <= ipv4.strm.dat;
          tcp.strm.sof <= pld_byte_cnt == 0;
          tcp.strm.eof <= (pld_byte_cnt == tcp.meta.pld_len - 1);
          tcp.strm.val <= 1;
        end
        rst_s : begin
          tcp.meta.val <= 1;
          tcp.strm.dat <= 0;
          tcp.strm.sof <= 0;
          tcp.strm.eof <= 0;
          tcp.strm.val <= 0;
          rst_reg      <= 1;
        end
      endcase
    end
  end
  //always_ff @ (posedge clk) if (rst) fsm_rst <= 1; else fsm_rst <= (tcp.strm.err || tcp.strm.eof);
  

endmodule : tcp_vlg_rx
