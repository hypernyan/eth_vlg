module bindfiles;
  bind mac_vlg_rx mac_vlg_rx_asrt p1 (.*);
endmodule : bindfiles