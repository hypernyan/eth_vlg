import ip_vlg_pkg::*;
import mac_vlg_pkg::*;
import eth_vlg_pkg::*;

interface ipv4
#( 
	parameter N = 1)
(
);

  logic      [7:0]  d;
  logic             v;
  logic             sof;
  logic             eof;
  logic             err;
  logic             busy;
  logic             done;
  logic             broadcast;
  length_t       payload_length;
  ipv4_hdr_t     ipv4_hdr;
  mac_hdr_t      mac_hdr;

  modport in_tx  (input  d, v, sof, eof, err, ipv4_hdr, mac_hdr, payload_length, broadcast, output busy, done); // used for transmitting ipv4 
  modport out_tx (output d, v, sof, eof, err, ipv4_hdr, mac_hdr, payload_length, broadcast, input  busy, done); // used for transmitting ipv4 

  modport in_rx  (input  d, v, sof, eof, err, ipv4_hdr, mac_hdr, payload_length); // used for receiving ipv4 
  modport out_rx (output d, v, sof, eof, err, ipv4_hdr, mac_hdr, payload_length); // used for receiving ipv4 
endinterface

module ip_vlg_top #(
  parameter int               N_TCP                = 1,
  parameter            [31:0] MTU                  = 1400,
  parameter [N_TCP-1:0][31:0] TCP_RETRANSMIT_TICKS = 1000000,
  parameter [N_TCP-1:0][31:0] TCP_RETRANSMIT_TRIES = 5,
  parameter [N_TCP-1:0][31:0] TCP_RAM_DEPTH        = 12,        
  parameter [N_TCP-1:0][31:0] TCP_PACKET_DEPTH     = 8,     
  parameter [N_TCP-1:0][31:0] TCP_WAIT_TICKS       = 100,
  parameter mac_addr_t        MAC_ADDR             = 0,
  parameter bit               DHCP_ENABLE          = 1,
  parameter int               DHCP_RETRIES         = 3
)
(
  input logic clk,
  input logic rst,
  mac.in      rx,
  mac.out     tx,
  input dev_t dev,
  input port_t [N_TCP-1:0] port,
  // Connects to ARP table
  output ipv4_t     ipv4_req,
  input  mac_addr_t mac_rsp,
  input  logic      arp_val,
  input  logic      arp_err,

  // Raw TCP
  input logic    [N_TCP-1:0]  [7:0] tcp_din,
  input logic    [N_TCP-1:0]        tcp_vin,
  output logic   [N_TCP-1:0]        tcp_cts,
  input logic    [N_TCP-1:0]        tcp_snd,

  output logic   [N_TCP-1:0]  [7:0] tcp_dout,
  output logic   [N_TCP-1:0]        tcp_vout,
  // TCP control [N_TCP-1:0]
  input  ipv4_t  [N_TCP-1:0]        rem_ipv4,
  input  port_t  [N_TCP-1:0]        rem_port,
  input  logic   [N_TCP-1:0]        connect, 
  output logic   [N_TCP-1:0]        connected,
  input  logic   [N_TCP-1:0]        listen,
  // Core status
  output logic   ready,
  output logic   error,
  // DHCP related
  input  ipv4_t  preferred_ipv4,
  output ipv4_t  assigned_ipv4,
  output logic   dhcp_success,
  output logic   dhcp_timeout
);

ipv4 ipv4_tx(.*);
ipv4 ipv4_rx(.*);

ipv4 icmp_ipv4_tx(.*);
ipv4 udp_ipv4_tx(.*);

udp udp_tx(.*);
udp udp_rx(.*);

ipv4_hdr_t [N_TCP+1:0] tx_ipv4_hdr_v;
mac_hdr_t  [N_TCP+1:0] tx_mac_hdr_v;
logic      [N_TCP+1:0] tx_mac_hdr_broadcast_v;

logic [N_TCP+1:0] act_ms;
logic rdy, avl;

wor   [N_TCP+1:0] ind;
logic [N_TCP+1:0] rst_fifo_vect;

ipv4_vlg ipv4_vlg_inst(
  .clk      (clk),
  .rst      (rst),
  .rst_fifo (rst_fifo),

  .mac_rx   (rx),
  .mac_tx   (tx),
  .dev      (dev),

  .rdy      (rdy),
  .avl      (avl),

  .ipv4_req (ipv4_req),
  .mac_rsp  (mac_rsp),
  .arp_val  (arp_val),
  .arp_err  (arp_err),
  .ipv4_tx  (ipv4_tx),
  .ipv4_rx  (ipv4_rx)
);

icmp_vlg icmp_vlg_inst (
  .clk  (clk),
  .rst  (rst),
  .rx   (ipv4_rx),
  .dev  (dev),
  .tx   (icmp_ipv4_tx)
);

udp_vlg udp_vlg_inst (
  .clk    (clk),
  .rst    (rst),
  .rx     (ipv4_rx),
  .tx     (udp_ipv4_tx),
  .udp_tx (udp_tx),
  .udp_rx (udp_rx),
  .dev    (dev)
);

dhcp_vlg #(
  .MAC_ADDR (MAC_ADDR),
  .ENABLE   (DHCP_ENABLE),
  .RETRIES  (DHCP_RETRIES)
) dhcp_vlg_inst (
  .clk (clk),
  .rst (rst),
  .rx  (udp_rx),
  .tx  (udp_tx),
 // .dev (dev),
  // Core status
  .ready (ready),
  .error (error),
  // DHCP related
  .preferred_ipv4 (preferred_ipv4),
  .assigned_ipv4  (assigned_ipv4),
  .dhcp_success   (dhcp_success),
  .dhcp_timeout   (dhcp_timeout)
);

logic [N_TCP-1:0][7:0] tcp_ipv4_tx_d;
logic [N_TCP-1:0]      tcp_ipv4_tx_v;

genvar i;

generate
  for (i = 0; i < N_TCP; i = i + 1) begin : gen_if
    ipv4 tcp_ipv4_tx(.*);
    ipv4 tcp_ipv4_rx(.*);
  end
endgenerate

generate 
  for (i = 0; i < N_TCP; i = i + 1) begin : gen_tcp
    tcp_vlg #(
      .MAX_PAYLOAD_LEN  (MTU - 120),
      .RETRANSMIT_TICKS (TCP_RETRANSMIT_TICKS[i]),
      .RETRANSMIT_TRIES (TCP_RETRANSMIT_TRIES[i]),
      .RAM_DEPTH        (TCP_RAM_DEPTH[i]),
      .PACKET_DEPTH     (TCP_PACKET_DEPTH[i]),
      .WAIT_TICKS       (TCP_WAIT_TICKS[i])
    ) tcp_vlg_inst (
      .clk       (clk),
      .rst       (rst),
      .dev       (dev),
      .port      (port[i]),
      .rx        (gen_if[i].tcp_ipv4_rx),
      .tx        (gen_if[i].tcp_ipv4_tx),
      .din       (tcp_din[i]),
      .vin       (tcp_vin[i]),
      .cts       (tcp_cts[i]),
      .snd       (tcp_snd[i]),

      .dout      (tcp_dout[i]),
      .vout      (tcp_vout[i]),

      .connected (connected[i]),
      .connect   (connect  [i]), 
      .listen    (listen   [i]),  
      .rem_ipv4  (rem_ipv4 [i]),
      .rem_port  (rem_port [i])
    );

    assign gen_if[i].tcp_ipv4_tx.done = ipv4_tx.eof && act_ms[i+2];
    assign gen_if[i].tcp_ipv4_tx.busy = ipv4_tx.busy;

    assign tcp_ipv4_tx_v[i] = gen_if[i].tcp_ipv4_tx.v;
    assign tcp_ipv4_tx_d[i] = gen_if[i].tcp_ipv4_tx.d;

    assign tx_ipv4_hdr_v[i+2]           = gen_if[i].tcp_ipv4_tx.ipv4_hdr;
    assign tx_mac_hdr_v [i+2]           = gen_if[i].tcp_ipv4_tx.mac_hdr;
    assign tx_mac_hdr_broadcast_v [i+2] = gen_if[i].tcp_ipv4_tx.broadcast;

    assign gen_if[i].tcp_ipv4_rx.d = ipv4_rx.d;
    assign gen_if[i].tcp_ipv4_rx.v = ipv4_rx.v;
    assign gen_if[i].tcp_ipv4_rx.sof = ipv4_rx.sof;
    assign gen_if[i].tcp_ipv4_rx.eof = ipv4_rx.eof;
    assign gen_if[i].tcp_ipv4_rx.err = ipv4_rx.err;
    assign gen_if[i].tcp_ipv4_rx.payload_length = ipv4_rx.payload_length;
    assign gen_if[i].tcp_ipv4_rx.ipv4_hdr = ipv4_rx.ipv4_hdr;
    assign gen_if[i].tcp_ipv4_rx.mac_hdr = ipv4_rx.mac_hdr;
  end
endgenerate

assign tx_ipv4_hdr_v[1]          = udp_ipv4_tx.ipv4_hdr;
assign tx_mac_hdr_v[1]           = udp_ipv4_tx.mac_hdr;
assign tx_mac_hdr_broadcast_v[1] = udp_ipv4_tx.broadcast;

assign tx_ipv4_hdr_v[0]          = icmp_ipv4_tx.ipv4_hdr;
assign tx_mac_hdr_v[0]           = icmp_ipv4_tx.mac_hdr;
assign tx_mac_hdr_broadcast_v[0] = icmp_ipv4_tx.broadcast;

generate
  for (i = 0; i < N_TCP + 2; i = i + 1) begin : gen_index
    assign ind = (act_ms[i] == 1'b1) ? i : 0;
    assign rst_fifo_vect[i] = (rst_fifo & act_ms[i]);
  end
endgenerate

assign icmp_ipv4_tx.done = ipv4_tx.eof && act_ms[0];
assign icmp_ipv4_tx.busy = ipv4_tx.busy;

assign ipv4_tx.ipv4_hdr = tx_ipv4_hdr_v[ind]; //
assign ipv4_tx.mac_hdr = tx_mac_hdr_v[ind]; //
assign ipv4_tx.broadcast = tx_mac_hdr_broadcast_v[ind]; //

buf_mng #(
  .W (8),
  .N (N_TCP + 2),
  .D ({{N_TCP{$clog2(MTU+1)}}, 32'h8, 32'd8}),
  .RWW (1)
)
buf_mng_inst (
  .clk (clk),
  .rst (rst),
  .rst_fifo (rst_fifo_vect), // flush fifo each sent IPv4 packet to avoid sending multiple packet's data if tcp or icmp continue to stream it.

  .v_i ({tcp_ipv4_tx_v[N_TCP-1:0], udp_ipv4_tx.v, icmp_ipv4_tx.v}),
  .d_i ({tcp_ipv4_tx_d[N_TCP-1:0], udp_ipv4_tx.d, icmp_ipv4_tx.d}),

  .v_o (ipv4_tx.v),
  .d_o (ipv4_tx.d),
  .eof (ipv4_tx.eof),
  .rdy (rdy),      // ipv4_tx is ready to accept data
  .avl (avl),      // data available to ipv4_tx
  .act_ms (act_ms) // tells which header to pass to ipv4_tx
);
endmodule

module ipv4_vlg (
  input logic clk,
  input logic rst,
  output logic rst_fifo,

  mac.in  mac_rx,
  mac.out mac_tx,
  input  dev_t dev,

  input  logic avl,
  output logic rdy,
// ARP request/response
  output ipv4_t    ipv4_req,
  input mac_addr_t mac_rsp,
  input logic      arp_val,
  input logic      arp_err,

  ipv4.in_tx  ipv4_tx,
  ipv4.out_rx ipv4_rx
);

mac_hdr_t mac_hdr;


ipv4_vlg_rx ipv4_vlg_rx_inst (
  .clk  (clk),
  .rst  (rst),
  .rx   (mac_rx),
  .ipv4 (ipv4_rx),
  .dev  (dev)
);


ipv4_vlg_tx ipv4_vlg_tx_inst (
  .clk  (clk),
  .rst  (rst),
  .rst_fifo (rst_fifo),
  .tx   (mac_tx),
  .ipv4 (ipv4_tx),
  .dev  (dev),
  .avl  (avl),
  .rdy  (rdy),

  .ipv4_req (ipv4_req),
  .mac_rsp  (mac_rsp),
  .arp_val  (arp_val),
  .arp_err  (arp_err)
);

endmodule : ipv4_vlg

module ipv4_vlg_rx #(
  parameter bit VERBOSE = 1
)
(
  input logic clk,
  input logic rst,
  mac.in      rx,
  ipv4.out_rx ipv4,
  input dev_t dev
);

// chsum

logic ipv4_v;
logic [7:0] ipv4_d;
logic ipv4_sof;
logic ipv4_eof;

assign ipv4_v = ipv4.v;
assign ipv4_d = ipv4.d;
assign ipv4_sof = ipv4.sof;
assign ipv4_eof = ipv4.eof;

logic [18:0] chsum;
logic [15:0] chsum_rec;
logic [15:0] chsum_calc;
logic [7:0]  chsum_hi;
logic [2:0]  chsum_carry;
logic        chsum_ctrl;
logic        chsum_ok;

assign chsum_carry = chsum[18:16];
assign chsum_calc  = chsum[15:0] + chsum_carry;

logic [15:0] byte_cnt;
logic fsm_rst, receiving, hdr_done;

logic [IPV4_HDR_LEN-1:0][7:0] hdr;

// Handle incoming packets, check for errors
logic [5:0] ihl_bytes;
always @ (posedge clk) begin
  if (fsm_rst || rst) begin
    receiving     <= 0;
    hdr_done      <= 0;
    chsum         <= 0;
    chsum_hi      <= 0;
    byte_cnt      <= 0;
    ipv4.d        <= 0;
    ipv4.sof      <= 0;
    ipv4.eof      <= 0;
    ipv4.ipv4_hdr <= 0;
  end
  else begin
    hdr[IPV4_HDR_LEN-1:1] <= hdr[IPV4_HDR_LEN-2:0];
    if (byte_cnt == IPV4_HDR_LEN-2) begin
      ipv4.ipv4_hdr[159:0] <= hdr[19:0];
      ipv4.payload_length <= hdr[17:16] - 20;
    end
    if (rx.sof && (rx.hdr.ethertype == eth_vlg_pkg::IPv4)) begin
      ihl_bytes <= {rx.d[3:0], 2'b00}; 
      receiving <= 1;
      $display("IPv4 RX");
    end
    if (receiving && (byte_cnt == (ihl_bytes - 1))) hdr_done <= 1;
    if (rx.v) begin
      if (byte_cnt[0]) chsum <= chsum + {chsum_hi, rx.d};
      if (!byte_cnt[0]) chsum_hi <= rx.d;
      if (receiving) byte_cnt <= byte_cnt + 1;
    end
    ipv4.d <= rx.d;
    ipv4.sof <= receiving && (byte_cnt == IPV4_HDR_LEN - 1);
    ipv4.eof <= hdr_done && (byte_cnt == ipv4.ipv4_hdr.length - 2);
  end
end

assign ipv4.v   = (hdr_done && (ipv4.ipv4_hdr.dst_ip == dev.ipv4_addr || ipv4.ipv4_hdr.dst_ip == IPV4_BROADCAST));
assign ipv4.err = rx.err;
assign fsm_rst  = (ipv4.eof || ipv4.err);
assign hdr[0] = rx.d;

// Calculate chsum
always @ (posedge clk) begin
  if (fsm_rst) begin
    chsum_ok <= 0;
  end
  else begin
    //if (chsum_ctrl && (chsum_calc == '1)) begin
    if (chsum_ctrl) begin
      chsum_ok <= 1;
    end
    else chsum_ok <= 0;
    if (chsum_ctrl && (chsum_calc != '1)) begin
      //if (fsm == ipv4_payload_s && byte_cnt == ipv4.ipv4_hdr.ihl*4) $display("IPv4 core: Bad header chsum.");
    end
  end
end

endmodule : ipv4_vlg_rx

module ipv4_vlg_tx #(
  parameter bit VERBOSE = 1
)
(
  input  logic  clk,
  input  logic  rst,
  output logic  rst_fifo,
  mac.out       tx,
  ipv4.in_tx    ipv4,
  input  dev_t  dev,
  input  logic  avl,
  output logic  rdy,
  // ARP table request/response
  output ipv4_t    ipv4_req,
  input mac_addr_t mac_rsp,
  input logic      arp_val,
  input logic      arp_err
);

localparam HDR_LEN = 20;

logic [7:0] ipv4_d;
logic ipv4_v;

assign ipv4_d = ipv4.d;
assign ipv4_v = ipv4.v;
logic ipv4_eof;
assign ipv4_eof = ipv4.eof;

logic fsm_rst;
logic hdr_done;

logic [HDR_LEN-1:0][7:0] hdr;
logic [HDR_LEN-1:0][7:0] hdr_calc;
logic [15:0] byte_cnt;


logic [15:0] chsum;
logic [18:0] chsum_carry;
logic [3:0] calc_byte_cnt;
logic calc;
logic calc_done;
logic [7:0] hdr_tx;

assign tx.hdr.src_mac_addr = dev.mac_addr;
assign arp_req_ipv4_addr = ipv4.ipv4_hdr.dst_ip;
assign rst_fifo = fsm_rst;

always @ (posedge clk) begin
  if (fsm_rst) begin
    calc           <= 0;
    hdr_calc       <= 0;
    chsum_carry    <= 0;
    calc_byte_cnt  <= 0;
    hdr_done       <= 0;
    calc_done      <= 0;
    byte_cnt       <= 0;
    rdy            <= 0;
    tx.v           <= 0;
    ipv4_req       <= 0;
    ipv4.busy      <= 0;
  end
  else begin
    if (avl && !ipv4.busy) begin // If data is available, latch the header for that data. !ipv4.busy to latch only once
      ipv4.busy         <= 1;
      hdr_calc[19]      <= {ipv4.ipv4_hdr.ver, ipv4.ipv4_hdr.ihl};
      hdr_calc[18]      <= ipv4.ipv4_hdr.qos;
      hdr_calc[17:16]   <= ipv4.ipv4_hdr.length;
      hdr_calc[15:14]   <= ipv4.ipv4_hdr.id;
      hdr_calc[13][7]   <= 0;
      hdr_calc[13][6]   <= ipv4.ipv4_hdr.df;
      hdr_calc[13][5]   <= ipv4.ipv4_hdr.mf;
      hdr_calc[13][4]   <= 0;
      hdr_calc[13][3:0] <= ipv4.ipv4_hdr.fo[11:8];
      hdr_calc[12]      <= ipv4.ipv4_hdr.fo[7:0];
      hdr_calc[11]      <= ipv4.ipv4_hdr.ttl;
      hdr_calc[10]      <= ipv4.ipv4_hdr.proto;
      hdr_calc[9:8]     <= 0;
      hdr_calc[7:4]     <= ipv4.ipv4_hdr.src_ip;
      hdr_calc[3:0]     <= ipv4.ipv4_hdr.dst_ip;
      calc <= 1; // Calculate chsum first
    end
    else if (calc) begin
      ipv4_req <= ipv4.ipv4_hdr.dst_ip; // Request MAC for destination IP
      calc_byte_cnt <= calc_byte_cnt + 1;
      chsum_carry <= chsum_carry + hdr_calc[1:0]; // Shift latched header and add up to chsum and carry
      hdr_calc[HDR_LEN-3:0] <= hdr_calc[HDR_LEN-1:2];
      if (calc_byte_cnt == 10) begin // Done with chsum
        calc_done <= 1; // Ready to readout data
        calc <= 0;
        hdr[19]      <= {ipv4.ipv4_hdr.ver, ipv4.ipv4_hdr.ihl};
        hdr[18]      <= ipv4.ipv4_hdr.qos;
        hdr[17:16]   <= ipv4.ipv4_hdr.length;
        hdr[15:14]   <= ipv4.ipv4_hdr.id;
        hdr[13][7]   <= 0;
        hdr[13][6]   <= ipv4.ipv4_hdr.df;
        hdr[13][5]   <= ipv4.ipv4_hdr.mf;
        hdr[13][4]   <= 0;
        hdr[13][3:0] <= ipv4.ipv4_hdr.fo[11:8];
        hdr[12]      <= ipv4.ipv4_hdr.fo[7:0];
        hdr[11]      <= ipv4.ipv4_hdr.ttl;
        hdr[10]      <= ipv4.ipv4_hdr.proto;
        hdr[9:8]     <= chsum;
        hdr[7:4]     <= ipv4.ipv4_hdr.src_ip;
        hdr[3:0]     <= ipv4.ipv4_hdr.dst_ip;
      end
    end
    if (calc_done && (arp_val || ipv4.broadcast)) begin // done calculating chsum, header completed now. ready to transmit when MAC from ARP table is valid
      tx.hdr.ethertype    <= eth_vlg_pkg::IPv4;
      tx.hdr.dst_mac_addr <= ipv4.broadcast ? '1 : mac_rsp; // acquire destination MAC from ARP table or assign it broadcast
      //tx.hdr.length       <= ipv4.ipv4_hdr.length + (ipv4.ipv4_hdr.ihl << 2);
      // if (byte_cnt == 0) $display ("<- srv: IPv4 to %d:%d:%d:%d.", hdr[3], hdr[2], hdr[1], hdr[0]);
      hdr[HDR_LEN-1:1] <= hdr[HDR_LEN-2:0];
      byte_cnt <= byte_cnt + 1;
      tx.sof <= (byte_cnt == 0);
      tx.v <= 1;
      if (byte_cnt == HDR_LEN-2) rdy <= 1;    // read out data from buffer. Buffer manager need 2 ticks to start output
      if (byte_cnt == HDR_LEN) hdr_done <= 1; // Done transmitting header, switch to buffer output
    end
  end
end

assign chsum = ~(chsum_carry[18:16] + chsum_carry[15:0]); // Calculate actual chsum
always @ (posedge clk) hdr_tx <= hdr[HDR_LEN-1];

assign tx.d = (hdr_done) ? ipv4.d : hdr_tx; // Switch data output between header and buffer's output
assign fsm_rst = (rst || ipv4.eof || arp_err);
assign tx.eof = ipv4.eof;
logic [7:0] txd;
logic txv;

assign txd = tx.d;
assign txv = tx.v;

endmodule : ipv4_vlg_tx
