import ipv4_vlg_pkg::*;
import mac_vlg_pkg::*;
import tcp_vlg_pkg::*;
import eth_vlg_pkg::*;

interface tcp;
  stream_t    strm;
  logic       rdy;   // data ready from to IPv4
  logic       req;   // data request for tx when done with header
  logic       ack;
  logic       done;
  tcp_meta_t  meta;

  modport in_rx  (input  strm, meta);
  modport out_rx (output strm, meta);
  modport in_tx  (input  strm, meta, rdy, output req, ack, done);
  modport out_tx (output strm, meta, rdy, input  req, ack, done);
endinterface : tcp

interface tcp_ctrl;
  logic  connect; 
  logic  listen;
  logic  connected;
  ipv4_t rem_ipv4;
  port_t rem_port;
  port_t loc_port;

  modport in  (input  connect, listen, rem_ipv4, rem_port, loc_port, output connected);
  modport out (output connect, listen, rem_ipv4, rem_port, loc_port, input  connected);
endinterface : tcp_ctrl

interface tcp_data;
  logic [7:0] dat; // data input
  logic       val; // data valid input
  logic       err; // error for rceive path only
  logic       cts; // transmission clear to send. user has 1 tick to deassert vin before data is lost
  logic       snd; // force sending all buffd data not waiting for TCP_WAIT_TICKS

  modport in_rx  (input  dat, val, err);
  modport out_rx (output dat, val, err);
  modport in_tx  (input  dat, val, snd, output cts);
  modport out_tx (output dat, val, snd, input  cts);
endinterface : tcp_data

interface rx_ctrl;
  logic     connected; // engine->rx_ctrl. connection established
  logic     flush;     // engine->rx_ctrl. request buffer flush
  logic     flushed;   // engine<-rx_ctrl. RAM flush successful
  tcb_t     tcb;       // engine->rx_ctrl. transmission control block
  stream_t  strm;      // engine->rx_ctrl. user data stream
  logic     init;      // engine->rx_ctrl. initialize loc_ack with tcb.loc_ack
  tcp_num_t loc_ack;   // engine<-rx_ctrl. current acknowledgement number (generated by rx control)
  logic     send_ack;  // force sending ack
  logic     ack_sent;

  modport in  (input  connected, flush, tcb, strm, init, ack_sent, output flushed, loc_ack, send_ack); 
  modport out (output connected, flush, tcb, strm, init, ack_sent, input  flushed, loc_ack, send_ack);
endinterface : rx_ctrl

interface tx_ctrl;
  logic     connected; // engine->tx_ctrl. connection established (generated by engine),
  logic     flush;     // engine->tx_ctrl. request buffer flush (generated by engine),
  logic     flushed;   // engine<-tx_ctrl. RAM was flushed (generated by buffer),
  tcb_t     tcb;       // engine->tx_ctrl. transmission control block wired from engine to rx and tx control,
  stream_t  strm;      // engine->tx_ctrl. user data stream,
  logic     init;      // engine->tx_ctrl. initialize loc_seq with tcb.loc_seq,
  tcp_num_t loc_seq;   // engine<-tx_ctrl. local sequence number,

  tcp_num_t pkt_seq;  // engine<-tx_ctrl. Transmitted packet's sequence number,

  length_t     len;       // engine<-tx_ctrl. packet's payload length,
  logic [31:0] cks;       // engine<-tx_ctrl. packet's payload checksum,
  logic        send;      // engine<-tx_ctrl. packet is ready for transmission (tx path only),
  logic        req;       // engine<-tx_ctrl. request strm (tx path only),
  logic        sent;      // engine<-tx_ctrl. tx is done,
  logic        force_dcn; // engine<-evt. force disconnect;
  modport in  (input  connected, flush, tcb, req, sent, init, output flushed, send, len, cks, strm, loc_seq, pkt_seq, force_dcn);
  modport out (output connected, flush, tcb, req, sent, init,  input flushed, send, len, cks, strm, loc_seq, pkt_seq, force_dcn);
endinterface : tx_ctrl
