import ipv4_vlg_pkg::*;
import mac_vlg_pkg::*;
import tcp_vlg_pkg::*;
import eth_vlg_pkg::*;

interface tcp;
  stream_t    strm;
  logic       rdy;  // data ready from to IPv4
  logic       req;  // data request for tx when done with header
  logic       acc;  // data accepted
  logic       done; // transmisssion finished
  tcp_meta_t  meta;

  modport in_rx  (input  strm, meta);
  modport out_rx (output strm, meta);
  modport in_tx  (input  strm, meta, rdy, output req, acc, done);
  modport out_tx (output strm, meta, rdy, input  req, acc, done);
endinterface : tcp

interface tcp_ctl;
  logic       connect; 
  logic       listen;
  tcp_stat_t  status;
  ipv4_t      rem_ipv4;
  port_t      rem_port;
  port_t      loc_port;

  modport in  (input  connect, listen, rem_ipv4, rem_port, loc_port, output status);
  modport out (output connect, listen, rem_ipv4, rem_port, loc_port, input  status);
endinterface : tcp_ctl

interface tcp_data;
  logic [7:0] dat; // data input
  logic       val; // data valid input
  logic       err; // error for rceive path only
  logic       cts; // transmission clear to send. user has 1 tick to deassert vin before data is lost
  logic       snd; // force sending all buffd data not waiting for TCP_WAIT_TICKS

  modport in_rx  (input  dat, val, err);
  modport out_rx (output dat, val, err);
  modport in_tx  (input  dat, val, snd, output cts);
  modport out_tx (output dat, val, snd, input  cts);
endinterface : tcp_data

interface rx_ctl;
  tcp_stat_t status; // engine->rx_ctl. connection established
  logic      flush;     // engine->rx_ctl. request buffer flush
  logic      flushed;   // engine<-rx_ctl. RAM flush successful
  tcb_t      tcb;       // engine->rx_ctl. transmission control block
  stream_t   strm;      // engine->rx_ctl. user data stream
  logic      init;      // engine->rx_ctl. initialize loc_ack with tcb.loc_ack
  tcp_num_t  loc_ack;   // engine<-rx_ctl. current acknowledgement number (generated by rx control)
  logic      send_ack;  // force sending ack
  logic      ack_sent;

  modport in  (input  status, flush, tcb, strm, init, ack_sent, output flushed, loc_ack, send_ack); 
  modport out (output status, flush, tcb, strm, init, ack_sent, input  flushed, loc_ack, send_ack);
endinterface : rx_ctl

interface tx_ctl;
  tcp_stat_t     status;    // engine->tx_ctl. connection established (generated by engine),
  logic          flush;     // engine->tx_ctl. request buffer flush (generated by engine),
  logic          flushed;   // engine<-tx_ctl. RAM was flushed (generated by buffer),
  tcb_t          tcb;       // engine->tx_ctl. transmission control block wired from engine to rx and tx control,
  stream_t       strm;      // engine->tx_ctl. user data stream,
  logic          init;      // engine->tx_ctl. initialize loc_seq with tcb.loc_seq,
  tcp_num_t      loc_seq;   // engine<-tx_ctl. local sequence number as in RAM's pointer
  logic          rst;       // engine->tx_ctl. reset transmission control
  tcp_pld_info_t pld_info;
  logic          send;      // engine<-tx_ctl. packet is ready for transmission (tx path only),
  logic          req;       // engine<-tx_ctl. request strm (tx path only),
  logic          sent;      // engine<-tx_ctl. tx is done,
  logic          force_dcn; // engine<-evt. force disconnect;
  modport in  (input  status, flush, tcb, req, sent, init, rst, output flushed, send, pld_info, strm, loc_seq, force_dcn);
  modport out (output status, flush, tcb, req, sent, init, rst,  input flushed, send, pld_info, strm, loc_seq, force_dcn);
endinterface : tx_ctl
