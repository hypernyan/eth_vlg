`define CLK_PERIOD 8
